library verilog;
use verilog.vl_types.all;
entity \OR\ is
    port(
        src0_i          : in     vl_logic;
        src1_i          : in     vl_logic;
        DataOut_o       : out    vl_logic
    );
end \OR\;
