library verilog;
use verilog.vl_types.all;
entity PC is
    port(
        clk             : in     vl_logic;
        new_PC          : in     vl_logic_vector(31 downto 0);
        PC_IFWrite      : in     vl_logic;
        rst_n           : in     vl_logic;
        PC_Addr         : out    vl_logic_vector(31 downto 0)
    );
end PC;
