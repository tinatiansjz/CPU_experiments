library verilog;
use verilog.vl_types.all;
entity IM_tb is
end IM_tb;
