module regfile(
  input clk,
  input rst_n,
  input Regwrite_i,

  input [4:0]wa_i, //rt or rd, write address
  input [4:0]ra0_i,//rs, read address 0 (Register number)
  input [4:0]ra1_i,//rt, read address 1 (Register number)
  input [31:0]wd_i,//write data
  output [31:0]rd0_o,  //rs, read data
  output [31:0]rd1_o   //rt, read data
  );
  reg [31:0] Regfile [31:0]; //31 31-bit register
  integer    i;
  always@(posedge clk or negedge rst_n)
  begin
    if (!rst_n)
      begin
        for (i = 1'b0; i < 32; i = i+1)
          Regfile[i] = 32'h0;
      end
    else
      begin
        if (Regwrite_i)
          Regfile[wa_i] = (!wa_i)? 32'h0 : wd_i;//only if the Regfile[wa_i] is not $zero
        
      end
  end
  //no other control inputs are needed. Read the content of the register anytime.
  assign rd0_o = Regfile[ra0_i];
  assign rd1_o = Regfile[ra1_i];
endmodule

