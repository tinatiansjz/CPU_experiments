library verilog;
use verilog.vl_types.all;
entity MIPS_tb is
end MIPS_tb;
